// CPU1.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU1 (
		output wire       buzzer_export,      //      buzzer.export
		input  wire       clk_clk,            //         clk.clk
		input  wire       key_1_export,       //       key_1.export
		input  wire       key_2_export,       //       key_2.export
		input  wire       key_3_export,       //       key_3.export
		output wire [9:0] leds_export,        //        leds.export
		input  wire       reset_reset_n,      //       reset.reset_n
		output wire [6:0] seven_seg_0_export, // seven_seg_0.export
		output wire [6:0] seven_seg_1_export, // seven_seg_1.export
		output wire [6:0] seven_seg_2_export, // seven_seg_2.export
		output wire [6:0] seven_seg_3_export, // seven_seg_3.export
		output wire [6:0] seven_seg_4_export, // seven_seg_4.export
		output wire [6:0] seven_seg_5_export, // seven_seg_5.export
		input  wire       sw_rst_export       //      sw_rst.export
	);

	wire  [31:0] cpu1_data_master_readdata;                                   // mm_interconnect_0:CPU1_data_master_readdata -> CPU1:d_readdata
	wire         cpu1_data_master_waitrequest;                                // mm_interconnect_0:CPU1_data_master_waitrequest -> CPU1:d_waitrequest
	wire         cpu1_data_master_debugaccess;                                // CPU1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU1_data_master_debugaccess
	wire  [13:0] cpu1_data_master_address;                                    // CPU1:d_address -> mm_interconnect_0:CPU1_data_master_address
	wire   [3:0] cpu1_data_master_byteenable;                                 // CPU1:d_byteenable -> mm_interconnect_0:CPU1_data_master_byteenable
	wire         cpu1_data_master_read;                                       // CPU1:d_read -> mm_interconnect_0:CPU1_data_master_read
	wire         cpu1_data_master_write;                                      // CPU1:d_write -> mm_interconnect_0:CPU1_data_master_write
	wire  [31:0] cpu1_data_master_writedata;                                  // CPU1:d_writedata -> mm_interconnect_0:CPU1_data_master_writedata
	wire  [31:0] cpu1_instruction_master_readdata;                            // mm_interconnect_0:CPU1_instruction_master_readdata -> CPU1:i_readdata
	wire         cpu1_instruction_master_waitrequest;                         // mm_interconnect_0:CPU1_instruction_master_waitrequest -> CPU1:i_waitrequest
	wire  [13:0] cpu1_instruction_master_address;                             // CPU1:i_address -> mm_interconnect_0:CPU1_instruction_master_address
	wire         cpu1_instruction_master_read;                                // CPU1:i_read -> mm_interconnect_0:CPU1_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_cpu1_debug_mem_slave_readdata;             // CPU1:debug_mem_slave_readdata -> mm_interconnect_0:CPU1_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu1_debug_mem_slave_waitrequest;          // CPU1:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU1_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu1_debug_mem_slave_debugaccess;          // mm_interconnect_0:CPU1_debug_mem_slave_debugaccess -> CPU1:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu1_debug_mem_slave_address;              // mm_interconnect_0:CPU1_debug_mem_slave_address -> CPU1:debug_mem_slave_address
	wire         mm_interconnect_0_cpu1_debug_mem_slave_read;                 // mm_interconnect_0:CPU1_debug_mem_slave_read -> CPU1:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu1_debug_mem_slave_byteenable;           // mm_interconnect_0:CPU1_debug_mem_slave_byteenable -> CPU1:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu1_debug_mem_slave_write;                // mm_interconnect_0:CPU1_debug_mem_slave_write -> CPU1:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu1_debug_mem_slave_writedata;            // mm_interconnect_0:CPU1_debug_mem_slave_writedata -> CPU1:debug_mem_slave_writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                        // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                          // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                           // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                             // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                         // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_key_1_s1_chipselect;                       // mm_interconnect_0:key_1_s1_chipselect -> key_1:chipselect
	wire  [31:0] mm_interconnect_0_key_1_s1_readdata;                         // key_1:readdata -> mm_interconnect_0:key_1_s1_readdata
	wire   [1:0] mm_interconnect_0_key_1_s1_address;                          // mm_interconnect_0:key_1_s1_address -> key_1:address
	wire         mm_interconnect_0_key_1_s1_write;                            // mm_interconnect_0:key_1_s1_write -> key_1:write_n
	wire  [31:0] mm_interconnect_0_key_1_s1_writedata;                        // mm_interconnect_0:key_1_s1_writedata -> key_1:writedata
	wire         mm_interconnect_0_key_2_s1_chipselect;                       // mm_interconnect_0:key_2_s1_chipselect -> key_2:chipselect
	wire  [31:0] mm_interconnect_0_key_2_s1_readdata;                         // key_2:readdata -> mm_interconnect_0:key_2_s1_readdata
	wire   [1:0] mm_interconnect_0_key_2_s1_address;                          // mm_interconnect_0:key_2_s1_address -> key_2:address
	wire         mm_interconnect_0_key_2_s1_write;                            // mm_interconnect_0:key_2_s1_write -> key_2:write_n
	wire  [31:0] mm_interconnect_0_key_2_s1_writedata;                        // mm_interconnect_0:key_2_s1_writedata -> key_2:writedata
	wire         mm_interconnect_0_key_3_s1_chipselect;                       // mm_interconnect_0:key_3_s1_chipselect -> key_3:chipselect
	wire  [31:0] mm_interconnect_0_key_3_s1_readdata;                         // key_3:readdata -> mm_interconnect_0:key_3_s1_readdata
	wire   [1:0] mm_interconnect_0_key_3_s1_address;                          // mm_interconnect_0:key_3_s1_address -> key_3:address
	wire         mm_interconnect_0_key_3_s1_write;                            // mm_interconnect_0:key_3_s1_write -> key_3:write_n
	wire  [31:0] mm_interconnect_0_key_3_s1_writedata;                        // mm_interconnect_0:key_3_s1_writedata -> key_3:writedata
	wire         mm_interconnect_0_seven_seg_0_s1_chipselect;                 // mm_interconnect_0:seven_seg_0_s1_chipselect -> seven_seg_0:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_readdata;                   // seven_seg_0:readdata -> mm_interconnect_0:seven_seg_0_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_0_s1_address;                    // mm_interconnect_0:seven_seg_0_s1_address -> seven_seg_0:address
	wire         mm_interconnect_0_seven_seg_0_s1_write;                      // mm_interconnect_0:seven_seg_0_s1_write -> seven_seg_0:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_0_s1_writedata;                  // mm_interconnect_0:seven_seg_0_s1_writedata -> seven_seg_0:writedata
	wire         mm_interconnect_0_seven_seg_1_s1_chipselect;                 // mm_interconnect_0:seven_seg_1_s1_chipselect -> seven_seg_1:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_readdata;                   // seven_seg_1:readdata -> mm_interconnect_0:seven_seg_1_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_1_s1_address;                    // mm_interconnect_0:seven_seg_1_s1_address -> seven_seg_1:address
	wire         mm_interconnect_0_seven_seg_1_s1_write;                      // mm_interconnect_0:seven_seg_1_s1_write -> seven_seg_1:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_1_s1_writedata;                  // mm_interconnect_0:seven_seg_1_s1_writedata -> seven_seg_1:writedata
	wire         mm_interconnect_0_seven_seg_2_s1_chipselect;                 // mm_interconnect_0:seven_seg_2_s1_chipselect -> seven_seg_2:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_readdata;                   // seven_seg_2:readdata -> mm_interconnect_0:seven_seg_2_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_2_s1_address;                    // mm_interconnect_0:seven_seg_2_s1_address -> seven_seg_2:address
	wire         mm_interconnect_0_seven_seg_2_s1_write;                      // mm_interconnect_0:seven_seg_2_s1_write -> seven_seg_2:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_2_s1_writedata;                  // mm_interconnect_0:seven_seg_2_s1_writedata -> seven_seg_2:writedata
	wire         mm_interconnect_0_seven_seg_3_s1_chipselect;                 // mm_interconnect_0:seven_seg_3_s1_chipselect -> seven_seg_3:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_readdata;                   // seven_seg_3:readdata -> mm_interconnect_0:seven_seg_3_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_3_s1_address;                    // mm_interconnect_0:seven_seg_3_s1_address -> seven_seg_3:address
	wire         mm_interconnect_0_seven_seg_3_s1_write;                      // mm_interconnect_0:seven_seg_3_s1_write -> seven_seg_3:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_3_s1_writedata;                  // mm_interconnect_0:seven_seg_3_s1_writedata -> seven_seg_3:writedata
	wire         mm_interconnect_0_seven_seg_4_s1_chipselect;                 // mm_interconnect_0:seven_seg_4_s1_chipselect -> seven_seg_4:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_readdata;                   // seven_seg_4:readdata -> mm_interconnect_0:seven_seg_4_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_4_s1_address;                    // mm_interconnect_0:seven_seg_4_s1_address -> seven_seg_4:address
	wire         mm_interconnect_0_seven_seg_4_s1_write;                      // mm_interconnect_0:seven_seg_4_s1_write -> seven_seg_4:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_4_s1_writedata;                  // mm_interconnect_0:seven_seg_4_s1_writedata -> seven_seg_4:writedata
	wire         mm_interconnect_0_seven_seg_5_s1_chipselect;                 // mm_interconnect_0:seven_seg_5_s1_chipselect -> seven_seg_5:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_5_s1_readdata;                   // seven_seg_5:readdata -> mm_interconnect_0:seven_seg_5_s1_readdata
	wire   [1:0] mm_interconnect_0_seven_seg_5_s1_address;                    // mm_interconnect_0:seven_seg_5_s1_address -> seven_seg_5:address
	wire         mm_interconnect_0_seven_seg_5_s1_write;                      // mm_interconnect_0:seven_seg_5_s1_write -> seven_seg_5:write_n
	wire  [31:0] mm_interconnect_0_seven_seg_5_s1_writedata;                  // mm_interconnect_0:seven_seg_5_s1_writedata -> seven_seg_5:writedata
	wire         mm_interconnect_0_ram_0_s1_chipselect;                       // mm_interconnect_0:ram_0_s1_chipselect -> ram_0:chipselect
	wire  [31:0] mm_interconnect_0_ram_0_s1_readdata;                         // ram_0:readdata -> mm_interconnect_0:ram_0_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_0_s1_address;                          // mm_interconnect_0:ram_0_s1_address -> ram_0:address
	wire   [3:0] mm_interconnect_0_ram_0_s1_byteenable;                       // mm_interconnect_0:ram_0_s1_byteenable -> ram_0:byteenable
	wire         mm_interconnect_0_ram_0_s1_write;                            // mm_interconnect_0:ram_0_s1_write -> ram_0:write
	wire  [31:0] mm_interconnect_0_ram_0_s1_writedata;                        // mm_interconnect_0:ram_0_s1_writedata -> ram_0:writedata
	wire         mm_interconnect_0_ram_0_s1_clken;                            // mm_interconnect_0:ram_0_s1_clken -> ram_0:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_buzzer_s1_chipselect;                      // mm_interconnect_0:buzzer_s1_chipselect -> buzzer:chipselect
	wire  [31:0] mm_interconnect_0_buzzer_s1_readdata;                        // buzzer:readdata -> mm_interconnect_0:buzzer_s1_readdata
	wire   [1:0] mm_interconnect_0_buzzer_s1_address;                         // mm_interconnect_0:buzzer_s1_address -> buzzer:address
	wire         mm_interconnect_0_buzzer_s1_write;                           // mm_interconnect_0:buzzer_s1_write -> buzzer:write_n
	wire  [31:0] mm_interconnect_0_buzzer_s1_writedata;                       // mm_interconnect_0:buzzer_s1_writedata -> buzzer:writedata
	wire  [31:0] mm_interconnect_0_sw_rst_s1_readdata;                        // sw_rst:readdata -> mm_interconnect_0:sw_rst_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_rst_s1_address;                         // mm_interconnect_0:sw_rst_s1_address -> sw_rst:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // key_1:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // key_2:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // key_3:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // timer_0:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu1_irq_irq;                                                // irq_mapper:sender_irq -> CPU1:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [CPU1:reset_n, buzzer:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, key_1:reset_n, key_2:reset_n, key_3:reset_n, leds:reset_n, mm_interconnect_0:CPU1_reset_reset_bridge_in_reset_reset, ram_0:reset, rst_translator:in_reset, seven_seg_0:reset_n, seven_seg_1:reset_n, seven_seg_2:reset_n, seven_seg_3:reset_n, seven_seg_4:reset_n, seven_seg_5:reset_n, sw_rst:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [CPU1:reset_req, ram_0:reset_req, rst_translator:reset_req_in]
	wire         cpu1_debug_reset_request_reset;                              // CPU1:debug_reset_request -> rst_controller:reset_in1

	CPU1_CPU1 cpu1 (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (cpu1_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu1_data_master_read),                              //                          .read
		.d_readdata                          (cpu1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu1_data_master_write),                             //                          .write
		.d_writedata                         (cpu1_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu1_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu1_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu1_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	CPU1_buzzer buzzer (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_buzzer_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_buzzer_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_buzzer_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_buzzer_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_buzzer_s1_readdata),   //                    .readdata
		.out_port   (buzzer_export)                           // external_connection.export
	);

	CPU1_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	CPU1_key_1 key_1 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_key_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_1_s1_readdata),   //                    .readdata
		.in_port    (key_1_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)               //                 irq.irq
	);

	CPU1_key_1 key_2 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_key_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_2_s1_readdata),   //                    .readdata
		.in_port    (key_2_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)               //                 irq.irq
	);

	CPU1_key_1 key_3 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_key_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_3_s1_readdata),   //                    .readdata
		.in_port    (key_3_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)               //                 irq.irq
	);

	CPU1_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	CPU1_ram_0 ram_0 (
		.clk        (clk_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_ram_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze     (1'b0)                                   // (terminated)
	);

	CPU1_seven_seg_0 seven_seg_0 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_0_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_0_export)                           // external_connection.export
	);

	CPU1_seven_seg_0 seven_seg_1 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_1_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_1_export)                           // external_connection.export
	);

	CPU1_seven_seg_0 seven_seg_2 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_2_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_2_export)                           // external_connection.export
	);

	CPU1_seven_seg_0 seven_seg_3 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_3_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_3_export)                           // external_connection.export
	);

	CPU1_seven_seg_0 seven_seg_4 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_4_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_4_export)                           // external_connection.export
	);

	CPU1_seven_seg_0 seven_seg_5 (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_seven_seg_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seven_seg_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seven_seg_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seven_seg_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seven_seg_5_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_5_export)                           // external_connection.export
	);

	CPU1_sw_rst sw_rst (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_sw_rst_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_rst_s1_readdata), //                    .readdata
		.in_port  (sw_rst_export)                         // external_connection.export
	);

	CPU1_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                 //   irq.irq
	);

	CPU1_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                        clk_0_clk.clk
		.CPU1_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                              // CPU1_reset_reset_bridge_in_reset.reset
		.CPU1_data_master_address                  (cpu1_data_master_address),                                    //                 CPU1_data_master.address
		.CPU1_data_master_waitrequest              (cpu1_data_master_waitrequest),                                //                                 .waitrequest
		.CPU1_data_master_byteenable               (cpu1_data_master_byteenable),                                 //                                 .byteenable
		.CPU1_data_master_read                     (cpu1_data_master_read),                                       //                                 .read
		.CPU1_data_master_readdata                 (cpu1_data_master_readdata),                                   //                                 .readdata
		.CPU1_data_master_write                    (cpu1_data_master_write),                                      //                                 .write
		.CPU1_data_master_writedata                (cpu1_data_master_writedata),                                  //                                 .writedata
		.CPU1_data_master_debugaccess              (cpu1_data_master_debugaccess),                                //                                 .debugaccess
		.CPU1_instruction_master_address           (cpu1_instruction_master_address),                             //          CPU1_instruction_master.address
		.CPU1_instruction_master_waitrequest       (cpu1_instruction_master_waitrequest),                         //                                 .waitrequest
		.CPU1_instruction_master_read              (cpu1_instruction_master_read),                                //                                 .read
		.CPU1_instruction_master_readdata          (cpu1_instruction_master_readdata),                            //                                 .readdata
		.buzzer_s1_address                         (mm_interconnect_0_buzzer_s1_address),                         //                        buzzer_s1.address
		.buzzer_s1_write                           (mm_interconnect_0_buzzer_s1_write),                           //                                 .write
		.buzzer_s1_readdata                        (mm_interconnect_0_buzzer_s1_readdata),                        //                                 .readdata
		.buzzer_s1_writedata                       (mm_interconnect_0_buzzer_s1_writedata),                       //                                 .writedata
		.buzzer_s1_chipselect                      (mm_interconnect_0_buzzer_s1_chipselect),                      //                                 .chipselect
		.CPU1_debug_mem_slave_address              (mm_interconnect_0_cpu1_debug_mem_slave_address),              //             CPU1_debug_mem_slave.address
		.CPU1_debug_mem_slave_write                (mm_interconnect_0_cpu1_debug_mem_slave_write),                //                                 .write
		.CPU1_debug_mem_slave_read                 (mm_interconnect_0_cpu1_debug_mem_slave_read),                 //                                 .read
		.CPU1_debug_mem_slave_readdata             (mm_interconnect_0_cpu1_debug_mem_slave_readdata),             //                                 .readdata
		.CPU1_debug_mem_slave_writedata            (mm_interconnect_0_cpu1_debug_mem_slave_writedata),            //                                 .writedata
		.CPU1_debug_mem_slave_byteenable           (mm_interconnect_0_cpu1_debug_mem_slave_byteenable),           //                                 .byteenable
		.CPU1_debug_mem_slave_waitrequest          (mm_interconnect_0_cpu1_debug_mem_slave_waitrequest),          //                                 .waitrequest
		.CPU1_debug_mem_slave_debugaccess          (mm_interconnect_0_cpu1_debug_mem_slave_debugaccess),          //                                 .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //    jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                 .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                 .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                 .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                 .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                 .chipselect
		.key_1_s1_address                          (mm_interconnect_0_key_1_s1_address),                          //                         key_1_s1.address
		.key_1_s1_write                            (mm_interconnect_0_key_1_s1_write),                            //                                 .write
		.key_1_s1_readdata                         (mm_interconnect_0_key_1_s1_readdata),                         //                                 .readdata
		.key_1_s1_writedata                        (mm_interconnect_0_key_1_s1_writedata),                        //                                 .writedata
		.key_1_s1_chipselect                       (mm_interconnect_0_key_1_s1_chipselect),                       //                                 .chipselect
		.key_2_s1_address                          (mm_interconnect_0_key_2_s1_address),                          //                         key_2_s1.address
		.key_2_s1_write                            (mm_interconnect_0_key_2_s1_write),                            //                                 .write
		.key_2_s1_readdata                         (mm_interconnect_0_key_2_s1_readdata),                         //                                 .readdata
		.key_2_s1_writedata                        (mm_interconnect_0_key_2_s1_writedata),                        //                                 .writedata
		.key_2_s1_chipselect                       (mm_interconnect_0_key_2_s1_chipselect),                       //                                 .chipselect
		.key_3_s1_address                          (mm_interconnect_0_key_3_s1_address),                          //                         key_3_s1.address
		.key_3_s1_write                            (mm_interconnect_0_key_3_s1_write),                            //                                 .write
		.key_3_s1_readdata                         (mm_interconnect_0_key_3_s1_readdata),                         //                                 .readdata
		.key_3_s1_writedata                        (mm_interconnect_0_key_3_s1_writedata),                        //                                 .writedata
		.key_3_s1_chipselect                       (mm_interconnect_0_key_3_s1_chipselect),                       //                                 .chipselect
		.leds_s1_address                           (mm_interconnect_0_leds_s1_address),                           //                          leds_s1.address
		.leds_s1_write                             (mm_interconnect_0_leds_s1_write),                             //                                 .write
		.leds_s1_readdata                          (mm_interconnect_0_leds_s1_readdata),                          //                                 .readdata
		.leds_s1_writedata                         (mm_interconnect_0_leds_s1_writedata),                         //                                 .writedata
		.leds_s1_chipselect                        (mm_interconnect_0_leds_s1_chipselect),                        //                                 .chipselect
		.ram_0_s1_address                          (mm_interconnect_0_ram_0_s1_address),                          //                         ram_0_s1.address
		.ram_0_s1_write                            (mm_interconnect_0_ram_0_s1_write),                            //                                 .write
		.ram_0_s1_readdata                         (mm_interconnect_0_ram_0_s1_readdata),                         //                                 .readdata
		.ram_0_s1_writedata                        (mm_interconnect_0_ram_0_s1_writedata),                        //                                 .writedata
		.ram_0_s1_byteenable                       (mm_interconnect_0_ram_0_s1_byteenable),                       //                                 .byteenable
		.ram_0_s1_chipselect                       (mm_interconnect_0_ram_0_s1_chipselect),                       //                                 .chipselect
		.ram_0_s1_clken                            (mm_interconnect_0_ram_0_s1_clken),                            //                                 .clken
		.seven_seg_0_s1_address                    (mm_interconnect_0_seven_seg_0_s1_address),                    //                   seven_seg_0_s1.address
		.seven_seg_0_s1_write                      (mm_interconnect_0_seven_seg_0_s1_write),                      //                                 .write
		.seven_seg_0_s1_readdata                   (mm_interconnect_0_seven_seg_0_s1_readdata),                   //                                 .readdata
		.seven_seg_0_s1_writedata                  (mm_interconnect_0_seven_seg_0_s1_writedata),                  //                                 .writedata
		.seven_seg_0_s1_chipselect                 (mm_interconnect_0_seven_seg_0_s1_chipselect),                 //                                 .chipselect
		.seven_seg_1_s1_address                    (mm_interconnect_0_seven_seg_1_s1_address),                    //                   seven_seg_1_s1.address
		.seven_seg_1_s1_write                      (mm_interconnect_0_seven_seg_1_s1_write),                      //                                 .write
		.seven_seg_1_s1_readdata                   (mm_interconnect_0_seven_seg_1_s1_readdata),                   //                                 .readdata
		.seven_seg_1_s1_writedata                  (mm_interconnect_0_seven_seg_1_s1_writedata),                  //                                 .writedata
		.seven_seg_1_s1_chipselect                 (mm_interconnect_0_seven_seg_1_s1_chipselect),                 //                                 .chipselect
		.seven_seg_2_s1_address                    (mm_interconnect_0_seven_seg_2_s1_address),                    //                   seven_seg_2_s1.address
		.seven_seg_2_s1_write                      (mm_interconnect_0_seven_seg_2_s1_write),                      //                                 .write
		.seven_seg_2_s1_readdata                   (mm_interconnect_0_seven_seg_2_s1_readdata),                   //                                 .readdata
		.seven_seg_2_s1_writedata                  (mm_interconnect_0_seven_seg_2_s1_writedata),                  //                                 .writedata
		.seven_seg_2_s1_chipselect                 (mm_interconnect_0_seven_seg_2_s1_chipselect),                 //                                 .chipselect
		.seven_seg_3_s1_address                    (mm_interconnect_0_seven_seg_3_s1_address),                    //                   seven_seg_3_s1.address
		.seven_seg_3_s1_write                      (mm_interconnect_0_seven_seg_3_s1_write),                      //                                 .write
		.seven_seg_3_s1_readdata                   (mm_interconnect_0_seven_seg_3_s1_readdata),                   //                                 .readdata
		.seven_seg_3_s1_writedata                  (mm_interconnect_0_seven_seg_3_s1_writedata),                  //                                 .writedata
		.seven_seg_3_s1_chipselect                 (mm_interconnect_0_seven_seg_3_s1_chipselect),                 //                                 .chipselect
		.seven_seg_4_s1_address                    (mm_interconnect_0_seven_seg_4_s1_address),                    //                   seven_seg_4_s1.address
		.seven_seg_4_s1_write                      (mm_interconnect_0_seven_seg_4_s1_write),                      //                                 .write
		.seven_seg_4_s1_readdata                   (mm_interconnect_0_seven_seg_4_s1_readdata),                   //                                 .readdata
		.seven_seg_4_s1_writedata                  (mm_interconnect_0_seven_seg_4_s1_writedata),                  //                                 .writedata
		.seven_seg_4_s1_chipselect                 (mm_interconnect_0_seven_seg_4_s1_chipselect),                 //                                 .chipselect
		.seven_seg_5_s1_address                    (mm_interconnect_0_seven_seg_5_s1_address),                    //                   seven_seg_5_s1.address
		.seven_seg_5_s1_write                      (mm_interconnect_0_seven_seg_5_s1_write),                      //                                 .write
		.seven_seg_5_s1_readdata                   (mm_interconnect_0_seven_seg_5_s1_readdata),                   //                                 .readdata
		.seven_seg_5_s1_writedata                  (mm_interconnect_0_seven_seg_5_s1_writedata),                  //                                 .writedata
		.seven_seg_5_s1_chipselect                 (mm_interconnect_0_seven_seg_5_s1_chipselect),                 //                                 .chipselect
		.sw_rst_s1_address                         (mm_interconnect_0_sw_rst_s1_address),                         //                        sw_rst_s1.address
		.sw_rst_s1_readdata                        (mm_interconnect_0_sw_rst_s1_readdata),                        //                                 .readdata
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                        //                       timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                          //                                 .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                       //                                 .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),                      //                                 .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect)                      //                                 .chipselect
	);

	CPU1_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu1_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu1_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
