// CPU1_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU1_tb (
	);

	wire        cpu1_inst_clk_bfm_clk_clk;           // CPU1_inst_clk_bfm:clk -> [CPU1_inst:clk_clk, CPU1_inst_reset_bfm:clk]
	wire        cpu1_inst_buzzer_export;             // CPU1_inst:buzzer_export -> CPU1_inst_buzzer_bfm:sig_export
	wire  [0:0] cpu1_inst_key_1_bfm_conduit_export;  // CPU1_inst_key_1_bfm:sig_export -> CPU1_inst:key_1_export
	wire  [0:0] cpu1_inst_key_2_bfm_conduit_export;  // CPU1_inst_key_2_bfm:sig_export -> CPU1_inst:key_2_export
	wire  [0:0] cpu1_inst_key_3_bfm_conduit_export;  // CPU1_inst_key_3_bfm:sig_export -> CPU1_inst:key_3_export
	wire  [9:0] cpu1_inst_leds_export;               // CPU1_inst:leds_export -> CPU1_inst_leds_bfm:sig_export
	wire  [6:0] cpu1_inst_seven_seg_0_export;        // CPU1_inst:seven_seg_0_export -> CPU1_inst_seven_seg_0_bfm:sig_export
	wire  [6:0] cpu1_inst_seven_seg_1_export;        // CPU1_inst:seven_seg_1_export -> CPU1_inst_seven_seg_1_bfm:sig_export
	wire  [6:0] cpu1_inst_seven_seg_2_export;        // CPU1_inst:seven_seg_2_export -> CPU1_inst_seven_seg_2_bfm:sig_export
	wire  [6:0] cpu1_inst_seven_seg_3_export;        // CPU1_inst:seven_seg_3_export -> CPU1_inst_seven_seg_3_bfm:sig_export
	wire  [6:0] cpu1_inst_seven_seg_4_export;        // CPU1_inst:seven_seg_4_export -> CPU1_inst_seven_seg_4_bfm:sig_export
	wire  [6:0] cpu1_inst_seven_seg_5_export;        // CPU1_inst:seven_seg_5_export -> CPU1_inst_seven_seg_5_bfm:sig_export
	wire  [0:0] cpu1_inst_sw_rst_bfm_conduit_export; // CPU1_inst_sw_rst_bfm:sig_export -> CPU1_inst:sw_rst_export
	wire        cpu1_inst_reset_bfm_reset_reset;     // CPU1_inst_reset_bfm:reset -> CPU1_inst:reset_reset_n

	CPU1 cpu1_inst (
		.buzzer_export      (cpu1_inst_buzzer_export),             //      buzzer.export
		.clk_clk            (cpu1_inst_clk_bfm_clk_clk),           //         clk.clk
		.key_1_export       (cpu1_inst_key_1_bfm_conduit_export),  //       key_1.export
		.key_2_export       (cpu1_inst_key_2_bfm_conduit_export),  //       key_2.export
		.key_3_export       (cpu1_inst_key_3_bfm_conduit_export),  //       key_3.export
		.leds_export        (cpu1_inst_leds_export),               //        leds.export
		.reset_reset_n      (cpu1_inst_reset_bfm_reset_reset),     //       reset.reset_n
		.seven_seg_0_export (cpu1_inst_seven_seg_0_export),        // seven_seg_0.export
		.seven_seg_1_export (cpu1_inst_seven_seg_1_export),        // seven_seg_1.export
		.seven_seg_2_export (cpu1_inst_seven_seg_2_export),        // seven_seg_2.export
		.seven_seg_3_export (cpu1_inst_seven_seg_3_export),        // seven_seg_3.export
		.seven_seg_4_export (cpu1_inst_seven_seg_4_export),        // seven_seg_4.export
		.seven_seg_5_export (cpu1_inst_seven_seg_5_export),        // seven_seg_5.export
		.sw_rst_export      (cpu1_inst_sw_rst_bfm_conduit_export)  //      sw_rst.export
	);

	altera_conduit_bfm cpu1_inst_buzzer_bfm (
		.sig_export (cpu1_inst_buzzer_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) cpu1_inst_clk_bfm (
		.clk (cpu1_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0002 cpu1_inst_key_1_bfm (
		.sig_export (cpu1_inst_key_1_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 cpu1_inst_key_2_bfm (
		.sig_export (cpu1_inst_key_2_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 cpu1_inst_key_3_bfm (
		.sig_export (cpu1_inst_key_3_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0003 cpu1_inst_leds_bfm (
		.sig_export (cpu1_inst_leds_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) cpu1_inst_reset_bfm (
		.reset (cpu1_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (cpu1_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0004 cpu1_inst_seven_seg_0_bfm (
		.sig_export (cpu1_inst_seven_seg_0_export)  // conduit.export
	);

	altera_conduit_bfm_0004 cpu1_inst_seven_seg_1_bfm (
		.sig_export (cpu1_inst_seven_seg_1_export)  // conduit.export
	);

	altera_conduit_bfm_0004 cpu1_inst_seven_seg_2_bfm (
		.sig_export (cpu1_inst_seven_seg_2_export)  // conduit.export
	);

	altera_conduit_bfm_0004 cpu1_inst_seven_seg_3_bfm (
		.sig_export (cpu1_inst_seven_seg_3_export)  // conduit.export
	);

	altera_conduit_bfm_0004 cpu1_inst_seven_seg_4_bfm (
		.sig_export (cpu1_inst_seven_seg_4_export)  // conduit.export
	);

	altera_conduit_bfm_0004 cpu1_inst_seven_seg_5_bfm (
		.sig_export (cpu1_inst_seven_seg_5_export)  // conduit.export
	);

	altera_conduit_bfm_0002 cpu1_inst_sw_rst_bfm (
		.sig_export (cpu1_inst_sw_rst_bfm_conduit_export)  // conduit.export
	);

endmodule
