// CPU1_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU1_tb (
	);

	wire        cpu1_inst_clk_bfm_clk_clk;       // CPU1_inst_clk_bfm:clk -> [CPU1_inst:clk_clk, CPU1_inst_reset_bfm:clk]
	wire  [1:0] cpu1_inst_leds_export;           // CPU1_inst:leds_export -> CPU1_inst_leds_bfm:sig_export
	wire        cpu1_inst_reset_bfm_reset_reset; // CPU1_inst_reset_bfm:reset -> CPU1_inst:reset_reset_n

	CPU1 cpu1_inst (
		.clk_clk            (cpu1_inst_clk_bfm_clk_clk),       //         clk.clk
		.key_1_export       (),                                //       key_1.export
		.key_2_export       (),                                //       key_2.export
		.key_3_export       (),                                //       key_3.export
		.leds_export        (cpu1_inst_leds_export),           //        leds.export
		.reset_reset_n      (cpu1_inst_reset_bfm_reset_reset), //       reset.reset_n
		.seven_seg_0_export (),                                // seven_seg_0.export
		.seven_seg_1_export (),                                // seven_seg_1.export
		.seven_seg_2_export (),                                // seven_seg_2.export
		.seven_seg_3_export (),                                // seven_seg_3.export
		.seven_seg_4_export (),                                // seven_seg_4.export
		.seven_seg_5_export ()                                 // seven_seg_5.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) cpu1_inst_clk_bfm (
		.clk (cpu1_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm cpu1_inst_leds_bfm (
		.sig_export (cpu1_inst_leds_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) cpu1_inst_reset_bfm (
		.reset (cpu1_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (cpu1_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
